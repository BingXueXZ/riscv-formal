//Need riscv formal interface